/*
PARAMETERS FOR PUF CONTROL MODULE
*/
parameter data_width = 32;
parameter addr_width = 32;
parameter puf_sig_length = 256;
parameter valid_byte_offset = 16;
parameter parity_bits_width = 48;