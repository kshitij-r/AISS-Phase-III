`define GPIO_IDATA 6'h5
`define GPIO_ODATA 6'h0

`define SYS_BUS_WAKEUP 24'b1000000
`define RST_Request 24'b1
`define Operation_Release_to_Host 24'b10000

`define IPID_N 0

`define CHIP_ID_ADDR 'h0
`define SECURE_COMMUNICATION_KEY_ADDR 'h1
`define LC_AUTHENTICATION_ID_ADDR_START 'h0


`define SCAN_KEY_WIDTH 64
`define SCAN_KEY_NUMBER 8